library verilog;
use verilog.vl_types.all;
entity Jiaotong_Lights_vlg_vec_tst is
end Jiaotong_Lights_vlg_vec_tst;
