`timescale 1ns/1ns
module tb_led();

//wire define
wire led_out ;
//reg define
reg key_in ;

//???????
initial key_in <= 1'b0;

//key_in:?????????????????
always #10 key_in <= {$random} % 2; /*?????????????0?1
??10ns???????*/

//------------- led_inst -------------
led led_inst
(
.key_in (key_in ), //input key_in

.led_out(led_out) //output led_out
);

endmodule
