library verilog;
use verilog.vl_types.all;
entity Jiaotong_lights_vlg_vec_tst is
end Jiaotong_lights_vlg_vec_tst;
