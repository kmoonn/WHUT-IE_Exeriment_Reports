library verilog;
use verilog.vl_types.all;
entity subway_vlg_vec_tst is
end subway_vlg_vec_tst;
